----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:42:55 08/09/2016 
-- Design Name: 
-- Module Name:    Transmitter_Core - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Transmitter_Core is
    Port ( Data_TX : in  STD_LOGIC_VECTOR (7 downto 0);
           Send : in  STD_LOGIC;
           TX : out  STD_LOGIC);
end Transmitter_Core;

architecture Behavioral of Transmitter_Core is

begin


end Behavioral;

